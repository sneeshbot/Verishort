module mod(a,b,c,d,e);
input a;
input b;
input c;
output d;
output e;
endmodule
