module mod(clock,reset,a);
	input clock;
	input reset;

	output a;
	assign a=1;
	endmodule
