module mod(a,b);
	input [11:0] a;
	output [11:0] b;
	assign b=a;
	endmodule
