module mod(_clock,_reset, a);
	input _clock;
	input _reset;
	output [3:0] a;
	assign a=15;
	endmodule
