module mod0(_clock,_reset,a,b);
	input _clock;
	input _reset;

	input a;
	output b;
	endmodule

module mod1(_clock,_reset,a,b);
	input _clock;
	input _reset;

	input a;
	output b;
	endmodule
