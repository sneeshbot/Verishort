module mod(clock,reset,a);
	input clock;
	input reset;

	output a;
	endmodule
