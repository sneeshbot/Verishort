module mod(_clock,_reset,a);
	input _clock;
	input _reset;

	output a;
	assign a=13'b0101010101011;
	endmodule
