module mod(a);
output a;
endmodule
