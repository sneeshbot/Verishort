module mod(clock,reset,a,b);
	input clock;
	input reset;

	input [20:0] a;
	output [30:0] b;
	endmodule
