module mod(_clock,_reset,a,b,c,d,e);
	input _clock;
	input _reset;
	input a;
	input b;
	input c;
	output d;
	output e;
	endmodule
