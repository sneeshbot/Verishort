module mod(_clock,_reset,a,b);
	input _clock;
	input _reset;

	input [20:0] a;
	output [30:0] b;
	endmodule
