module mod(a, b);
input a;
output b;
endmodule
