module m(b,c,x,y);
	output [1:0] b;
	output c;
	output x;
	output [2:0] y;
	
	wire [1:0]a;
	wire d;
	wire e;
	wire [2:0]f;
	
	assign b=a;
	assign c=d;
	assign x=e;
	assign y=f;
	endmodule
