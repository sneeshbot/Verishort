module mod(clock,reset,a);
	input clock;
	input reset;

	output a;
	assign a=0'b0101010101011;
	endmodule
