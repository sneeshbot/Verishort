module mod(clock,reset, a);
	input clock;
	input reset;
	output [3:0] a;
	a=15;
	endmodule
