module mod(a,b);
	input [20:0] a;
	output [30:0] b;
	endmodule
