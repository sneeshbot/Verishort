module mod(_clock,_reset,a);
	input _clock;
	input _reset;

	output a;
	endmodule
