module mod(a);
	output a;
	assign a=0'b0101010101011;
	endmodule
