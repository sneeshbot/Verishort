module a();
	wire [10:0]b;
	assign b = 1;
	endmodule
