module mod0(a,b);
input a;
output b;
endmodule

module mod1(a,b);
input a;
output b;
endmodule
