module mod(clock,reset,a, b);
	input clock;
	input reset;

	input a;
	output b;
	endmodule
