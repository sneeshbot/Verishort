module mod(a,b,c);
	input [9:0] a;
	input b;
	output c;
	assign c=a;
	endmodule
