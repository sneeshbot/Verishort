module mod(clock,reset,a,b,c,d,e);
	input clock;
	input reset;
	input a;
	input b;
	input c;
	output d;
	output e;
	endmodule
