module mod(_clock,_reset,a, b);
	input _clock;
	input _reset;

	input a;
	output b;
	endmodule
