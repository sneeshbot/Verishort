module mod(a);
	output [3:0] a;
	a=15;
	endmodule
