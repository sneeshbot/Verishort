module mod(a)
	output a;
	assign a=1;
	endmodule;
