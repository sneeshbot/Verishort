module mod0(clock,reset,a,b);
	input clock;
	input reset;

	input a;
	output b;
	endmodule

module mod1(clock,reset,a,b);
	input clock;
	input reset;

	input a;
	output b;
	endmodule
